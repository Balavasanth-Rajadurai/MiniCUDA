
`default_nettype none
`timescale 1ns/1ns

module controller #(
    parameter ADDR_BITS = 8,
    parameter DATA_BITS = 16,
    parameter NUM_CONSUMERS = 4,
    parameter NUM_CHANNELS = 1,
    parameter WRITE_ENABLE = 1
)(
    input  wire clk,
    input  wire reset,

    input  wire [NUM_CONSUMERS-1:0]                      consumer_read_valid,
    input  wire [ADDR_BITS-1:0]                          consumer_read_address  [NUM_CONSUMERS-1:0],
    output reg  [NUM_CONSUMERS-1:0]                      consumer_read_ready,
    output reg  [DATA_BITS-1:0]                          consumer_read_data     [NUM_CONSUMERS-1:0],

    input  wire [NUM_CONSUMERS-1:0]                      consumer_write_valid,
    input  wire [ADDR_BITS-1:0]                          consumer_write_address [NUM_CONSUMERS-1:0],
    input  wire [DATA_BITS-1:0]                          consumer_write_data    [NUM_CONSUMERS-1:0],
    output reg  [NUM_CONSUMERS-1:0]                      consumer_write_ready,

    output reg  [NUM_CHANNELS-1:0]                       mem_read_valid,
    output reg  [ADDR_BITS-1:0]                          mem_read_address       [NUM_CHANNELS-1:0],
    input  wire [NUM_CHANNELS-1:0]                       mem_read_ready,
    input  wire [DATA_BITS-1:0]                          mem_read_data          [NUM_CHANNELS-1:0],

    output reg  [NUM_CHANNELS-1:0]                       mem_write_valid,
    output reg  [ADDR_BITS-1:0]                          mem_write_address      [NUM_CHANNELS-1:0],
    output reg  [DATA_BITS-1:0]                          mem_write_data         [NUM_CHANNELS-1:0],
    input  wire [NUM_CHANNELS-1:0]                       mem_write_ready
);

    localparam IDLE           = 3'b000,
               READ_WAITING   = 3'b010,
               WRITE_WAITING  = 3'b011,
               READ_RELAYING  = 3'b100,
               WRITE_RELAYING = 3'b101;

    reg [2:0] controller_state [NUM_CHANNELS-1:0];
    reg [$clog2(NUM_CONSUMERS)-1:0] current_consumer [NUM_CHANNELS-1:0];
    reg [NUM_CONSUMERS-1:0] channel_serving_consumer [NUM_CHANNELS-1:0];

    integer i, j;

    always @(posedge clk) begin
        if (reset) begin
            for (i = 0; i < NUM_CHANNELS; i++) begin
                controller_state[i] <= IDLE;
                mem_read_valid[i]   <= 0;
                mem_write_valid[i]  <= 0;
                mem_read_address[i] <= 0;
                mem_write_address[i]<= 0;
                mem_write_data[i]   <= 0;
                current_consumer[i] <= 0;

                for (j = 0; j < NUM_CONSUMERS; j++) begin
                    channel_serving_consumer[i][j] <= 0;
                    consumer_read_ready[j]         <= 0;
                    consumer_write_ready[j]        <= 0;
                    consumer_read_data[j]          <= 0;
                end
            end
        end else begin
            for (i = 0; i < NUM_CHANNELS; i++) begin
                case (controller_state[i])
                    IDLE: begin : inner_loop
                        for (j = 0; j < NUM_CONSUMERS; j++) begin
                            if (consumer_read_valid[j] && !channel_serving_consumer[i][j]) begin
                                channel_serving_consumer[i][j] <= 1;
                                current_consumer[i]            <= j;
                                mem_read_valid[i]              <= 1;
                                mem_read_address[i]            <= consumer_read_address[j];
                                controller_state[i]            <= READ_WAITING;
                                disable inner_loop;
                            end else if (consumer_write_valid[j] && !channel_serving_consumer[i][j]) begin
                                channel_serving_consumer[i][j] <= 1;
                                current_consumer[i]            <= j;
                                mem_write_valid[i]             <= 1;
                                mem_write_address[i]           <= consumer_write_address[j];
                                mem_write_data[i]              <= consumer_write_data[j];
                                controller_state[i]            <= WRITE_WAITING;
                                disable inner_loop;
                            end
                        end
                    end

                    READ_WAITING: begin
                        if (mem_read_ready[i]) begin
                            mem_read_valid[i]                          <= 0;
                            consumer_read_ready[current_consumer[i]]   <= 1;
                            consumer_read_data[current_consumer[i]]    <= mem_read_data[i];
                            controller_state[i]                        <= READ_RELAYING;
                        end
                    end

                    WRITE_WAITING: begin
                        if (mem_write_ready[i]) begin
                            mem_write_valid[i]                         <= 0;
                            consumer_write_ready[current_consumer[i]]  <= 1;
                            controller_state[i]                        <= WRITE_RELAYING;
                        end
                    end

                    READ_RELAYING: begin
                        if (!consumer_read_valid[current_consumer[i]]) begin
                            channel_serving_consumer[i][current_consumer[i]] <= 0;
                            consumer_read_ready[current_consumer[i]]         <= 0;
                            controller_state[i]                              <= IDLE;
                        end
                    end

                    WRITE_RELAYING: begin
                        if (!consumer_write_valid[current_consumer[i]]) begin
                            channel_serving_consumer[i][current_consumer[i]] <= 0;
                            consumer_write_ready[current_consumer[i]]        <= 0;
                            controller_state[i]                              <= IDLE;
                        end
                    end
                endcase
            end
        end
    end

endmodule

